v {xschem version=3.4.8RC file_version=1.2}
G {}
K {}
V {}
S {}
E {}
N -30 -70 -30 -50 {lab=vnmic}
N -30 -70 20 -70 {lab=vnmic}
N 80 -70 110 -70 {lab=vn1}
N 170 -70 210 -70 {lab=vn2}
N -30 10 -30 50 {lab=GND}
N 300 -210 330 -210 {lab=#net1}
N 300 -210 300 -70 {lab=#net1}
N 280 -70 320 -70 {lab=#net1}
N 270 -70 280 -70 {lab=#net1}
N 300 -150 330 -150 {lab=#net1}
N 430 -50 430 -10 {lab=GND}
N 390 -150 420 -150 {lab=vout}
N 390 -210 430 -210 {lab=vout}
N 420 -150 430 -150 {lab=vout}
N 430 -210 430 -120 {lab=vout}
N 430 -60 430 -50 {lab=GND}
N 360 20 360 40 {lab=GND}
N 360 40 360 70 {lab=GND}
N 590 -40 590 0 {lab=GND}
N 360 -100 380 -100 {lab=vcm}
N 360 -100 360 -40 {lab=vcm}
N 320 -70 370 -70 {lab=#net1}
N 370 -80 380 -80 {lab=#net1}
N 370 -80 370 -70 {lab=#net1}
N 430 -120 500 -120 {lab=vout}
N 500 -120 510 -120 {lab=vout}
N 510 -120 510 -90 {lab=vout}
N 540 -100 590 -100 {lab=vout}
N 540 -100 540 -90 {lab=vout}
N 510 -90 540 -90 {lab=vout}
N 430 -60 450 -60 {lab=GND}
C {vsource.sym} -30 -20 0 0 {name=Vmic value="0 AC 1" savecurrent=false}
C {capa.sym} 140 -70 3 0 {name=C1
m=1
value=4.7u
footprint=1206
device="ceramic capacitor"}
C {gnd.sym} 430 -10 0 0 {name=l1 lab=GND}
C {res.sym} 50 -70 3 0 {name=R1
value=380
footprint=1206
device=resistor
m=1}
C {res.sym} 240 -70 3 0 {name=R2
value=4.7k
footprint=1206
device=resistor
m=1}
C {gnd.sym} -30 50 0 0 {name=l2 lab=GND}
C {capa.sym} 360 -210 3 0 {name=C2
m=1
value=27u
footprint=1206
device="ceramic capacitor"}
C {res.sym} 360 -150 3 0 {name=R3
value=300k
footprint=1206
device=resistor
m=1}
C {vsource.sym} 360 -10 0 0 {name=V2 value=1.5 savecurrent=false}
C {capa.sym} 590 -70 0 0 {name=C3
m=1
value=4.7u
footprint=1206
device="ceramic capacitor"}
C {gnd.sym} 360 70 0 0 {name=l3 lab=GND}
C {gnd.sym} 590 0 0 0 {name=l4 lab=GND}
C {simulator_commands_shown.sym} 920 -410 0 0 {name=COMMANDS
simulator=ngspice
only_toplevel=false 
value="
.CONTROL

OP
save all
write mydesign.raw
set appendwrite
AC DEC 100 0.1 10e6
write mydesign.raw
MEAS AC gain_db MAX vdb(vout) FROM=0.1 TO=10e6
LET vm3db=gain_db-3.0
print vm3db
.ENDC
"}
C {lab_wire.sym} 13.37347800263035 -70 0 0 {name=p1 sig_type=std_logic lab=vnmic}
C {lab_wire.sym} 90 -70 1 0 {name=p2 sig_type=std_logic lab=vn1}
C {lab_wire.sym} 180 -70 1 0 {name=p3 sig_type=std_logic lab=vn2}
C {lab_wire.sym} 360 -40 0 0 {name=p4 sig_type=std_logic lab=vcm}
C {lab_wire.sym} 510 -90 1 0 {name=p5 sig_type=std_logic lab=vout}
C {opamp.sym} 620 100 0 0 {name=x1}
